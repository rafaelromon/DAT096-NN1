
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY LINE_BUFF_tb IS
	GENERIC
	(
		INPUT_WIDTH     : INTEGER := 9;
		INPUT_HEIGHT    : INTEGER := 9;
		INPUT_CHANNELS  : INTEGER := 1;
		FILTERS         : INTEGER := 1;
		KERNEL_HEIGHT   : INTEGER := 3;
		KERNEL_WIDTH    : INTEGER := 3;
		KERNEL_CHANNELS : INTEGER := 1;
		INTEGER_SIZE    : INTEGER := 8
	);
END LINE_BUFF_tb;

ARCHITECTURE LINE_BUFF_tb_arch OF LINE_BUFF_tb IS

	SIGNAL clk_tb     : STD_LOGIC := '1';
	SIGNAL reset_p_tb : STD_LOGIC := '0';
	SIGNAL start_tb   : STD_LOGIC := '0';
	SIGNAL input_tb   : STD_LOGIC_VECTOR((INPUT_WIDTH * INPUT_HEIGHT * INTEGER_SIZE) - 1 DOWNTO 0);
	SIGNAL busy_tb    : STD_LOGIC;
	SIGNAL done_tb    : STD_LOGIC;
	SIGNAL output_tb  : STD_LOGIC_VECTOR((KERNEL_HEIGHT * KERNEL_WIDTH * INTEGER_SIZE) - 1 DOWNTO 0);

	COMPONENT LINE_BUFF
		GENERIC
		(
			INPUT_WIDTH    : INTEGER := 128;
			INPUT_HEIGHT   : INTEGER := 128;
			INPUT_CHANNELS : INTEGER := 8;
			KERNEL_WIDTH   : INTEGER := 1;
			KERNEL_HEIGHT  : INTEGER := 1;
			STRIDE         : INTEGER := 1;
			INTEGER_SIZE   : INTEGER := 8
		);
		PORT
		(
			clk     : IN  STD_LOGIC;
			reset_p : IN  STD_LOGIC;
			start   : IN  STD_LOGIC;
			move    : IN  STD_LOGIC;
			input   : IN  STD_LOGIC_VECTOR((INPUT_WIDTH * INPUT_HEIGHT * INTEGER_SIZE) - 1 DOWNTO 0);
			busy    : OUT STD_LOGIC;
			done    : OUT STD_LOGIC;
			output  : OUT STD_LOGIC_VECTOR((KERNEL_HEIGHT * KERNEL_WIDTH * INTEGER_SIZE) - 1 DOWNTO 0)
		);
	END COMPONENT LINE_BUFF;
BEGIN

	LINE_BUFF_i : LINE_BUFF
	GENERIC
	MAP (
	INPUT_WIDTH    => INPUT_WIDTH,
	INPUT_HEIGHT   => INPUT_HEIGHT,
	INPUT_CHANNELS => INPUT_CHANNELS,
	KERNEL_WIDTH   => KERNEL_WIDTH,
	KERNEL_HEIGHT  => KERNEL_HEIGHT,
	STRIDE         => 1,
	INTEGER_SIZE   => INTEGER_SIZE
	)
	PORT MAP
	(
		clk     => clk_tb,
		reset_p => reset_p_tb,
		start   => start_tb,
		move    => '1',
		input   => input_tb,
		busy    => busy_tb,
		done    => done_tb,
		output  => output_tb
	);

	clk_tb <= NOT clk_tb AFTER 10 ns;

	PROCESS IS
	BEGIN

		reset_p_tb <= '1';
		WAIT FOR 20ns;
		reset_p_tb <= '0';
		WAIT FOR 20ns;
		input_tb <= "000001001100000011010110001100010111000001111101010101010000111011001111001110101000010110110100111011110010111111101111101000010001100110100000110111110010111000100001011011110010101100010101001011011101100000110000101001000010101010111101000111000000010101111001100100010000100111100101001011110000000111010111010111010001101111001001100100000011001011000000101010100111000111001100101001010010001111011010001111011111011101100110110101011111111011101001111010010010101011110110100110011110101100010000100101001000000111011110101001010001011100101011110011111001011011110100111100111010001110000111011001111000000010001101110011101100110011111111";
		--input_tb <= "101101110010010100011000111000100111101010000001101111101111010101111010";
		start_tb <= '1';
		WAIT FOR 20ns;
		start_tb <= '0';
		WAIT FOR 10000ms;

	END PROCESS;

END LINE_BUFF_tb_arch;
