
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY PWConv_tb is
  generic (
    INPUT_WIDTH     : INTEGER := 9;
    INPUT_HEIGHT    : INTEGER := 9;
    INPUT_CHANNELS  : INTEGER := 1;
    FILTERS         : INTEGER := 1;
    KERNEL_HEIGHT   : INTEGER := 3;
    KERNEL_WIDTH    : INTEGER := 3;
    KERNEL_CHANNELS : INTEGER := 1;
    IN_SIZE         : INTEGER := 8;
    OUT_SIZE        : INTEGER := 32
  );
END PWConv_tb;

ARCHITECTURE PWConv_tb_arch OF PWConv_tb IS

signal clk_tb           : STD_LOGIC := '1';
signal reset_p_tb       : STD_LOGIC := '0';
signal enable_tb        : STD_LOGIC := '0';
signal input_tb         : STD_LOGIC_VECTOR((INPUT_WIDTH*INPUT_HEIGHT*IN_SIZE) - 1 DOWNTO 0);
signal filter_values_tb : STD_LOGIC_VECTOR ((FILTERS*KERNEL_HEIGHT*KERNEL_WIDTH*KERNEL_CHANNELS*IN_SIZE) - 1 DOWNTO 0);
signal bias_values_tb   : STD_LOGIC_VECTOR(OUT_SIZE - 1 DOWNTO 0);
signal busy_tb          : STD_LOGIC;
signal done_tb          : STD_LOGIC;
signal output_tb        : STD_LOGIC_VECTOR(OUT_SIZE - 1 DOWNTO 0);

component PWConv
generic (
  INPUT_WIDTH     : INTEGER := 128;
  INPUT_HEIGHT    : INTEGER := 128;
  INPUT_CHANNELS  : INTEGER := 8;
  FILTERS         : INTEGER := 32;
  KERNEL_HEIGHT   : INTEGER := 1;
  KERNEL_WIDTH    : INTEGER := 1;
  KERNEL_CHANNELS : INTEGER := 8;
  IN_SIZE         : INTEGER := 8;
  OUT_SIZE        : INTEGER := 32
);
port (
  clk           : IN  STD_LOGIC;
  reset_p       : IN  STD_LOGIC;
  enable        : IN  STD_LOGIC;
  input         : IN  STD_LOGIC_VECTOR((INPUT_WIDTH*INPUT_HEIGHT*IN_SIZE) - 1 DOWNTO 0);
  filter_values : IN  STD_LOGIC_VECTOR ((FILTERS*KERNEL_HEIGHT*KERNEL_WIDTH*KERNEL_CHANNELS*IN_SIZE) - 1 DOWNTO 0);
  bias_values   : IN  STD_LOGIC_VECTOR(FILTERS*OUT_SIZE - 1 DOWNTO 0);
  busy          : OUT STD_LOGIC;
  done          : OUT STD_LOGIC;
  output        : OUT STD_LOGIC_VECTOR(OUT_SIZE - 1 DOWNTO 0)
);
end component PWConv;

BEGIN

PWConv_i : PWConv
  generic map (
  INPUT_WIDTH     => INPUT_WIDTH,
  INPUT_HEIGHT    => INPUT_HEIGHT,
  INPUT_CHANNELS  => INPUT_CHANNELS,
  FILTERS         => FILTERS,
  KERNEL_HEIGHT   => KERNEL_HEIGHT,
  KERNEL_WIDTH    => KERNEL_WIDTH,
  KERNEL_CHANNELS => KERNEL_CHANNELS,
  IN_SIZE         => IN_SIZE,
  OUT_SIZE        => OUT_SIZE
  )
  port map (
  clk           => clk_tb,
  reset_p       => reset_p_tb,
  enable        => enable_tb,
  input         => input_tb,
  filter_values => filter_values_tb,
  bias_values   => bias_values_tb,
  busy          => busy_tb,
  done          => done_tb,
  output        => output_tb
  );


	clk_tb <= NOT clk_tb AFTER 10 ns;

	PROCESS IS
	BEGIN

		reset_p_tb <= '1';
		WAIT FOR 20ns;
		reset_p_tb <= '0';
		WAIT FOR 20ns;
		input_tb <= "000001001100000011010110001100010111000001111101010101010000111011001111001110101000010110110100111011110010111111101111101000010001100110100000110111110010111000100001011011110010101100010101001011011101100000110000101001000010101010111101000111000000010101111001100100010000100111100101001011110000000111010111010111010001101111001001100100000011001011000000101010100111000111001100101001010010001111011010001111011111011101100110110101011111111011101001111010010010101011110110100110011110101100010000100101001000000111011110101001010001011100101011110011111001011011110100111100111010001110000111011001111000000010001101110011101100110011111111";
        filter_values_tb <= "101101110010010100011000111000100111101010000001101111101111010101111010";
		bias_values_tb <= "10000101101101001110111100101111";
		enable_tb <= '1';
		WAIT FOR 20ns;
		enable_tb <= '0';
		WAIT FOR 10000ms;

	END PROCESS;

END PWConv_tb_arch;
