-----------------------------------------------------
-- Title: TOP_LEVEL.vhdl
-- Author: Rafael Rom�n/NN-1
-- DAT096 - spring 2021
-----------------------------------------------------
-- Description:
-- This entity dictates the top level
-- architecture of the entire system
-- TODO:
-- * implement BRAM controller
-- * better implement user button
-----------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY TOP_LEVEL IS
	PORT
	(
		SYSCLK_P     : IN STD_LOGIC;
		CPU_RESET    : IN STD_LOGIC;
		GPIO_SW_N    : IN STD_LOGIC;
		USB_UART_TX  : OUT STD_LOGIC;
		USB_UART_RTS : OUT STD_LOGIC
	);
END TOP_LEVEL;

ARCHITECTURE TOP_LEVEL_arch OF TOP_LEVEL IS

	TYPE states IS (Idle, LoadImage, ProcessImage, SendResult);
	SIGNAL state_machine : states := Idle;
	SIGNAL reset_signal: STD_LOGIC := '0';

	SIGNAL cnn_start : STD_LOGIC := '0';
	SIGNAL loaded_image : STD_LOGIC_VECTOR(16383 DOWNTO 0);
	SIGNAL cnn_finished : STD_LOGIC;
	SIGNAL cnn_result : STD_LOGIC_VECTOR(5 DOWNTO 0);

	COMPONENT CNN IS
		PORT
		(
			clk       : IN std_logic;
			reset_p   : IN std_logic;
			start     : IN std_logic;
			image     : IN std_logic_vector(16383 DOWNTO 0);
			finished  : OUT std_logic;
			result    : OUT std_logic_vector(5 DOWNTO 0)
		);
	END COMPONENT CNN;

	SIGNAL TX_DV : STD_LOGIC := '0';
	SIGNAL TX_Byte : STD_LOGIC_vector(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL TX_Done : STD_LOGIC;

	COMPONENT UART_TX IS
		PORT
		(
			clk        : IN STD_LOGIC;
			TX_DV      : IN STD_LOGIC;
			TX_Byte    : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			TX_Active  : OUT STD_LOGIC;
			TX_Serial  : OUT STD_LOGIC;
			TX_Done    : OUT STD_LOGIC
		);
	END COMPONENT UART_TX;

BEGIN
	CNN_comp : CNN -- Instantiate CNN transmitter
	PORT MAP
	(
		clk       => SYSCLK_P,
		reset_p   => reset_signal,
		start     => cnn_start,
		image     => loaded_image,
		finished  => cnn_finished,
		result    => cnn_result
	);

	UART_TX_comp : UART_TX -- Instantiate UART transmitter
	PORT MAP
	(
		clk        => SYSCLK_P,
		TX_DV      => TX_DV,
		TX_Byte    => TX_Byte,
		TX_Active  => USB_UART_RTS,
		TX_Serial  => USB_UART_TX,
		TX_Done    => TX_Done
	);

	-- Purpose: Control state machine
	TOP_LEVEL_process : PROCESS (SYSCLK_P, CPU_RESET)
	BEGIN
	    IF CPU_RESET = '1' THEN
           state_machine <= Idle;

		ELSIF RISING_EDGE(SYSCLK_P) THEN
			CASE state_machine IS
				WHEN Idle =>

					IF GPIO_SW_N = '0' THEN -- TODO this will cause problems once moved into the board
						reset_signal <= '0';
						state_machine <= LoadImage;
					ELSE
						reset_signal <= '1';
					END IF;

				WHEN LoadImage =>
					-- TODO this does nothing at the moment
					loaded_image <= (OTHERS => '0');
					state_machine <= ProcessImage;

				WHEN ProcessImage =>

					IF cnn_finished = '1' THEN
						cnn_start <= '0';
					    state_machine <= SendResult;
					ELSE
						cnn_start <= '1';
                    END IF;

				WHEN SendResult =>

					IF TX_DONE = '1' THEN
						TX_DV <= '0';
						state_machine <= Idle;
					ELSE
						TX_DV <= '1';
						TX_BYTE <= cnn_result;
					END IF;

			END CASE;
		END IF;
	END PROCESS TOP_LEVEL_process;
END TOP_LEVEL_arch;
