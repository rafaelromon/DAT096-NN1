-----------------------------------------------------
-- Title: PWConv.vhdl
-- Author: Rafael Romon/NN-1
-- DAT096 - spring 2021
-----------------------------------------------------
-- Description:
-- TODO:
-- Channels are not implemented
-----------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY PWConv IS

END PWConv;

ARCHITECTURE PWConv_arch OF PWConv IS
BEGIN
END PWConv_arch;
